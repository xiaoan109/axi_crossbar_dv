package axi_test_pkg;
  import uvm_pkg::*;
  // `include "uvm_macros.svh"

  import axi_stimulus_pkg::*;
  import axi_env_pkg::*;

  `include "axi_base_test.sv"
endpackage
