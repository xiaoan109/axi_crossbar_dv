`timescale 1ns / 10ps

module tb_top ();

  import uvm_pkg::*;
  import axi_globals_pkg::*;
  import axi_test_pkg::*;

  bit aclk;
  bit aresetn;
  bit srst;

  axi_if #(
      .AXI_DATA_W(AXI_DATA_W),
      .AXI_ADDR_W(AXI_ADDR_W),
      .AXI_ID_W  (AXI_ID_W),
      .AXI_USER_W(AXI_USER_W)
  ) mst[3:0] (
      .*
  );

  axi_if #(
      .AXI_DATA_W(AXI_DATA_W),
      .AXI_ADDR_W(AXI_ADDR_W),
      .AXI_ID_W  (AXI_ID_W),
      .AXI_USER_W(AXI_USER_W)
  ) slv[3:0] (
      .*
  );


  axicb_crossbar_top #(
      .AXI_ADDR_W     (AXI_ADDR_W),
      .AXI_ID_W       (AXI_ID_W),
      .AXI_DATA_W     (AXI_DATA_W),
      .MST_PIPELINE   (0),
      .SLV_PIPELINE   (0),
      .AXI_SIGNALING  (1),                // AXI Full
      .USER_SUPPORT   (1),
      .AXI_AUSER_W    (AXI_USER_W),
      .AXI_WUSER_W    (AXI_USER_W),
      .AXI_BUSER_W    (AXI_USER_W),
      .AXI_RUSER_W    (AXI_USER_W),
      .MST0_ID_MASK   (MST0_ID_MASK),
      .MST1_ID_MASK   (MST1_ID_MASK),
      .MST2_ID_MASK   (MST2_ID_MASK),
      .MST3_ID_MASK   (MST3_ID_MASK),
      .SLV0_START_ADDR(SLV0_START_ADDR),
      .SLV0_END_ADDR  (SLV0_END_ADDR),
      .SLV1_START_ADDR(SLV1_START_ADDR),
      .SLV1_END_ADDR  (SLV1_END_ADDR),
      .SLV2_START_ADDR(SLV2_START_ADDR),
      .SLV2_END_ADDR  (SLV2_END_ADDR),
      .SLV3_START_ADDR(SLV3_START_ADDR),
      .SLV3_END_ADDR  (SLV3_END_ADDR)
  ) dut (
      .aclk         (aclk),
      .aresetn      (aresetn),
      .srst         (srst),
      .slv0_aclk    (aclk),
      .slv0_aresetn (aresetn),
      .slv0_srst    (srst),
      .slv0_awvalid (mst[0].awvalid),
      .slv0_awready (mst[0].awready),
      .slv0_awaddr  (mst[0].awaddr),
      .slv0_awlen   (mst[0].awlen),
      .slv0_awsize  (mst[0].awsize),
      .slv0_awburst (mst[0].awburst),
      .slv0_awlock  (mst[0].awlock),
      .slv0_awcache (mst[0].awcache),
      .slv0_awprot  (mst[0].awprot),
      .slv0_awqos   (mst[0].awqos),
      .slv0_awregion(mst[0].awregion),
      .slv0_awid    (mst[0].awid),
      .slv0_awuser  (mst[0].awuser),
      .slv0_wvalid  (mst[0].wvalid),
      .slv0_wready  (mst[0].wready),
      .slv0_wlast   (mst[0].wlast),
      .slv0_wdata   (mst[0].wdata),
      .slv0_wstrb   (mst[0].wstrb),
      .slv0_wuser   (mst[0].wuser),
      .slv0_bvalid  (mst[0].bvalid),
      .slv0_bready  (mst[0].bready),
      .slv0_bid     (mst[0].bid),
      .slv0_bresp   (mst[0].bresp),
      .slv0_buser   (mst[0].buser),
      .slv0_arvalid (mst[0].arvalid),
      .slv0_arready (mst[0].arready),
      .slv0_araddr  (mst[0].araddr),
      .slv0_arlen   (mst[0].arlen),
      .slv0_arsize  (mst[0].arsize),
      .slv0_arburst (mst[0].arburst),
      .slv0_arlock  (mst[0].arlock),
      .slv0_arcache (mst[0].arcache),
      .slv0_arprot  (mst[0].arprot),
      .slv0_arqos   (mst[0].arqos),
      .slv0_arregion(mst[0].arregion),
      .slv0_arid    (mst[0].arid),
      .slv0_aruser  (mst[0].aruser),
      .slv0_rvalid  (mst[0].rvalid),
      .slv0_rready  (mst[0].rready),
      .slv0_rid     (mst[0].rid),
      .slv0_rresp   (mst[0].rresp),
      .slv0_rdata   (mst[0].rdata),
      .slv0_rlast   (mst[0].rlast),
      .slv0_ruser   (mst[0].ruser),
      .slv1_aclk    (aclk),
      .slv1_aresetn (aresetn),
      .slv1_srst    (srst),
      .slv1_awvalid (mst[1].awvalid),
      .slv1_awready (mst[1].awready),
      .slv1_awaddr  (mst[1].awaddr),
      .slv1_awlen   (mst[1].awlen),
      .slv1_awsize  (mst[1].awsize),
      .slv1_awburst (mst[1].awburst),
      .slv1_awlock  (mst[1].awlock),
      .slv1_awcache (mst[1].awcache),
      .slv1_awprot  (mst[1].awprot),
      .slv1_awqos   (mst[1].awqos),
      .slv1_awregion(mst[1].awregion),
      .slv1_awid    (mst[1].awid),
      .slv1_awuser  (mst[1].awuser),
      .slv1_wvalid  (mst[1].wvalid),
      .slv1_wready  (mst[1].wready),
      .slv1_wlast   (mst[1].wlast),
      .slv1_wdata   (mst[1].wdata),
      .slv1_wstrb   (mst[1].wstrb),
      .slv1_wuser   (mst[1].wuser),
      .slv1_bvalid  (mst[1].bvalid),
      .slv1_bready  (mst[1].bready),
      .slv1_bid     (mst[1].bid),
      .slv1_bresp   (mst[1].bresp),
      .slv1_buser   (mst[1].buser),
      .slv1_arvalid (mst[1].arvalid),
      .slv1_arready (mst[1].arready),
      .slv1_araddr  (mst[1].araddr),
      .slv1_arlen   (mst[1].arlen),
      .slv1_arsize  (mst[1].arsize),
      .slv1_arburst (mst[1].arburst),
      .slv1_arlock  (mst[1].arlock),
      .slv1_arcache (mst[1].arcache),
      .slv1_arprot  (mst[1].arprot),
      .slv1_arqos   (mst[1].arqos),
      .slv1_arregion(mst[1].arregion),
      .slv1_arid    (mst[1].arid),
      .slv1_aruser  (mst[1].aruser),
      .slv1_rvalid  (mst[1].rvalid),
      .slv1_rready  (mst[1].rready),
      .slv1_rid     (mst[1].rid),
      .slv1_rresp   (mst[1].rresp),
      .slv1_rdata   (mst[1].rdata),
      .slv1_rlast   (mst[1].rlast),
      .slv1_ruser   (mst[1].ruser),
      .slv2_aclk    (aclk),
      .slv2_aresetn (aresetn),
      .slv2_srst    (srst),
      .slv2_awvalid (mst[2].awvalid),
      .slv2_awready (mst[2].awready),
      .slv2_awaddr  (mst[2].awaddr),
      .slv2_awlen   (mst[2].awlen),
      .slv2_awsize  (mst[2].awsize),
      .slv2_awburst (mst[2].awburst),
      .slv2_awlock  (mst[2].awlock),
      .slv2_awcache (mst[2].awcache),
      .slv2_awprot  (mst[2].awprot),
      .slv2_awqos   (mst[2].awqos),
      .slv2_awregion(mst[2].awregion),
      .slv2_awid    (mst[2].awid),
      .slv2_awuser  (mst[2].awuser),
      .slv2_wvalid  (mst[2].wvalid),
      .slv2_wready  (mst[2].wready),
      .slv2_wlast   (mst[2].wlast),
      .slv2_wdata   (mst[2].wdata),
      .slv2_wstrb   (mst[2].wstrb),
      .slv2_wuser   (mst[2].wuser),
      .slv2_bvalid  (mst[2].bvalid),
      .slv2_bready  (mst[2].bready),
      .slv2_bid     (mst[2].bid),
      .slv2_bresp   (mst[2].bresp),
      .slv2_buser   (mst[2].buser),
      .slv2_arvalid (mst[2].arvalid),
      .slv2_arready (mst[2].arready),
      .slv2_araddr  (mst[2].araddr),
      .slv2_arlen   (mst[2].arlen),
      .slv2_arsize  (mst[2].arsize),
      .slv2_arburst (mst[2].arburst),
      .slv2_arlock  (mst[2].arlock),
      .slv2_arcache (mst[2].arcache),
      .slv2_arprot  (mst[2].arprot),
      .slv2_arqos   (mst[2].arqos),
      .slv2_arregion(mst[2].arregion),
      .slv2_arid    (mst[2].arid),
      .slv2_aruser  (mst[2].aruser),
      .slv2_rvalid  (mst[2].rvalid),
      .slv2_rready  (mst[2].rready),
      .slv2_rid     (mst[2].rid),
      .slv2_rresp   (mst[2].rresp),
      .slv2_rdata   (mst[2].rdata),
      .slv2_rlast   (mst[2].rlast),
      .slv2_ruser   (mst[2].ruser),
      .slv3_aclk    (aclk),
      .slv3_aresetn (aresetn),
      .slv3_srst    (srst),
      .slv3_awvalid (mst[3].awvalid),
      .slv3_awready (mst[3].awready),
      .slv3_awaddr  (mst[3].awaddr),
      .slv3_awlen   (mst[3].awlen),
      .slv3_awsize  (mst[3].awsize),
      .slv3_awburst (mst[3].awburst),
      .slv3_awlock  (mst[3].awlock),
      .slv3_awcache (mst[3].awcache),
      .slv3_awprot  (mst[3].awprot),
      .slv3_awqos   (mst[3].awqos),
      .slv3_awregion(mst[3].awregion),
      .slv3_awid    (mst[3].awid),
      .slv3_awuser  (mst[3].awuser),
      .slv3_wvalid  (mst[3].wvalid),
      .slv3_wready  (mst[3].wready),
      .slv3_wlast   (mst[3].wlast),
      .slv3_wdata   (mst[3].wdata),
      .slv3_wstrb   (mst[3].wstrb),
      .slv3_wuser   (mst[3].wuser),
      .slv3_bvalid  (mst[3].bvalid),
      .slv3_bready  (mst[3].bready),
      .slv3_bid     (mst[3].bid),
      .slv3_bresp   (mst[3].bresp),
      .slv3_buser   (mst[3].buser),
      .slv3_arvalid (mst[3].arvalid),
      .slv3_arready (mst[3].arready),
      .slv3_araddr  (mst[3].araddr),
      .slv3_arlen   (mst[3].arlen),
      .slv3_arsize  (mst[3].arsize),
      .slv3_arburst (mst[3].arburst),
      .slv3_arlock  (mst[3].arlock),
      .slv3_arcache (mst[3].arcache),
      .slv3_arprot  (mst[3].arprot),
      .slv3_arqos   (mst[3].arqos),
      .slv3_arregion(mst[3].arregion),
      .slv3_arid    (mst[3].arid),
      .slv3_aruser  (mst[3].aruser),
      .slv3_rvalid  (mst[3].rvalid),
      .slv3_rready  (mst[3].rready),
      .slv3_rid     (mst[3].rid),
      .slv3_rresp   (mst[3].rresp),
      .slv3_rdata   (mst[3].rdata),
      .slv3_rlast   (mst[3].rlast),
      .slv3_ruser   (mst[3].ruser),
      .mst0_aclk    (aclk),
      .mst0_aresetn (aresetn),
      .mst0_srst    (srst),
      .mst0_awvalid (slv[0].awvalid),
      .mst0_awready (slv[0].awready),
      .mst0_awaddr  (slv[0].awaddr),
      .mst0_awlen   (slv[0].awlen),
      .mst0_awsize  (slv[0].awsize),
      .mst0_awburst (slv[0].awburst),
      .mst0_awlock  (slv[0].awlock),
      .mst0_awcache (slv[0].awcache),
      .mst0_awprot  (slv[0].awprot),
      .mst0_awqos   (slv[0].awqos),
      .mst0_awregion(slv[0].awregion),
      .mst0_awid    (slv[0].awid),
      .mst0_awuser  (slv[0].awuser),
      .mst0_wvalid  (slv[0].wvalid),
      .mst0_wready  (slv[0].wready),
      .mst0_wlast   (slv[0].wlast),
      .mst0_wdata   (slv[0].wdata),
      .mst0_wstrb   (slv[0].wstrb),
      .mst0_wuser   (slv[0].wuser),
      .mst0_bvalid  (slv[0].bvalid),
      .mst0_bready  (slv[0].bready),
      .mst0_bid     (slv[0].bid),
      .mst0_bresp   (slv[0].bresp),
      .mst0_buser   (slv[0].buser),
      .mst0_arvalid (slv[0].arvalid),
      .mst0_arready (slv[0].arready),
      .mst0_araddr  (slv[0].araddr),
      .mst0_arlen   (slv[0].arlen),
      .mst0_arsize  (slv[0].arsize),
      .mst0_arburst (slv[0].arburst),
      .mst0_arlock  (slv[0].arlock),
      .mst0_arcache (slv[0].arcache),
      .mst0_arprot  (slv[0].arprot),
      .mst0_arqos   (slv[0].arqos),
      .mst0_arregion(slv[0].arregion),
      .mst0_arid    (slv[0].arid),
      .mst0_aruser  (slv[0].aruser),
      .mst0_rvalid  (slv[0].rvalid),
      .mst0_rready  (slv[0].rready),
      .mst0_rid     (slv[0].rid),
      .mst0_rresp   (slv[0].rresp),
      .mst0_rdata   (slv[0].rdata),
      .mst0_rlast   (slv[0].rlast),
      .mst0_ruser   (slv[0].ruser),
      .mst1_aclk    (aclk),
      .mst1_aresetn (aresetn),
      .mst1_srst    (srst),
      .mst1_awvalid (slv[1].awvalid),
      .mst1_awready (slv[1].awready),
      .mst1_awaddr  (slv[1].awaddr),
      .mst1_awlen   (slv[1].awlen),
      .mst1_awsize  (slv[1].awsize),
      .mst1_awburst (slv[1].awburst),
      .mst1_awlock  (slv[1].awlock),
      .mst1_awcache (slv[1].awcache),
      .mst1_awprot  (slv[1].awprot),
      .mst1_awqos   (slv[1].awqos),
      .mst1_awregion(slv[1].awregion),
      .mst1_awid    (slv[1].awid),
      .mst1_awuser  (slv[1].awuser),
      .mst1_wvalid  (slv[1].wvalid),
      .mst1_wready  (slv[1].wready),
      .mst1_wlast   (slv[1].wlast),
      .mst1_wdata   (slv[1].wdata),
      .mst1_wstrb   (slv[1].wstrb),
      .mst1_wuser   (slv[1].wuser),
      .mst1_bvalid  (slv[1].bvalid),
      .mst1_bready  (slv[1].bready),
      .mst1_bid     (slv[1].bid),
      .mst1_bresp   (slv[1].bresp),
      .mst1_buser   (slv[1].buser),
      .mst1_arvalid (slv[1].arvalid),
      .mst1_arready (slv[1].arready),
      .mst1_araddr  (slv[1].araddr),
      .mst1_arlen   (slv[1].arlen),
      .mst1_arsize  (slv[1].arsize),
      .mst1_arburst (slv[1].arburst),
      .mst1_arlock  (slv[1].arlock),
      .mst1_arcache (slv[1].arcache),
      .mst1_arprot  (slv[1].arprot),
      .mst1_arqos   (slv[1].arqos),
      .mst1_arregion(slv[1].arregion),
      .mst1_arid    (slv[1].arid),
      .mst1_aruser  (slv[1].aruser),
      .mst1_rvalid  (slv[1].rvalid),
      .mst1_rready  (slv[1].rready),
      .mst1_rid     (slv[1].rid),
      .mst1_rresp   (slv[1].rresp),
      .mst1_rdata   (slv[1].rdata),
      .mst1_rlast   (slv[1].rlast),
      .mst1_ruser   (slv[1].ruser),
      .mst2_aclk    (aclk),
      .mst2_aresetn (aresetn),
      .mst2_srst    (srst),
      .mst2_awvalid (slv[2].awvalid),
      .mst2_awready (slv[2].awready),
      .mst2_awaddr  (slv[2].awaddr),
      .mst2_awlen   (slv[2].awlen),
      .mst2_awsize  (slv[2].awsize),
      .mst2_awburst (slv[2].awburst),
      .mst2_awlock  (slv[2].awlock),
      .mst2_awcache (slv[2].awcache),
      .mst2_awprot  (slv[2].awprot),
      .mst2_awqos   (slv[2].awqos),
      .mst2_awregion(slv[2].awregion),
      .mst2_awid    (slv[2].awid),
      .mst2_awuser  (slv[2].awuser),
      .mst2_wvalid  (slv[2].wvalid),
      .mst2_wready  (slv[2].wready),
      .mst2_wlast   (slv[2].wlast),
      .mst2_wdata   (slv[2].wdata),
      .mst2_wstrb   (slv[2].wstrb),
      .mst2_wuser   (slv[2].wuser),
      .mst2_bvalid  (slv[2].bvalid),
      .mst2_bready  (slv[2].bready),
      .mst2_bid     (slv[2].bid),
      .mst2_bresp   (slv[2].bresp),
      .mst2_buser   (slv[2].buser),
      .mst2_arvalid (slv[2].arvalid),
      .mst2_arready (slv[2].arready),
      .mst2_araddr  (slv[2].araddr),
      .mst2_arlen   (slv[2].arlen),
      .mst2_arsize  (slv[2].arsize),
      .mst2_arburst (slv[2].arburst),
      .mst2_arlock  (slv[2].arlock),
      .mst2_arcache (slv[2].arcache),
      .mst2_arprot  (slv[2].arprot),
      .mst2_arqos   (slv[2].arqos),
      .mst2_arregion(slv[2].arregion),
      .mst2_arid    (slv[2].arid),
      .mst2_aruser  (slv[2].aruser),
      .mst2_rvalid  (slv[2].rvalid),
      .mst2_rready  (slv[2].rready),
      .mst2_rid     (slv[2].rid),
      .mst2_rresp   (slv[2].rresp),
      .mst2_rdata   (slv[2].rdata),
      .mst2_rlast   (slv[2].rlast),
      .mst2_ruser   (slv[2].ruser),
      .mst3_aclk    (aclk),
      .mst3_aresetn (aresetn),
      .mst3_srst    (srst),
      .mst3_awvalid (slv[3].awvalid),
      .mst3_awready (slv[3].awready),
      .mst3_awaddr  (slv[3].awaddr),
      .mst3_awlen   (slv[3].awlen),
      .mst3_awsize  (slv[3].awsize),
      .mst3_awburst (slv[3].awburst),
      .mst3_awlock  (slv[3].awlock),
      .mst3_awcache (slv[3].awcache),
      .mst3_awprot  (slv[3].awprot),
      .mst3_awqos   (slv[3].awqos),
      .mst3_awregion(slv[3].awregion),
      .mst3_awid    (slv[3].awid),
      .mst3_awuser  (slv[3].awuser),
      .mst3_wvalid  (slv[3].wvalid),
      .mst3_wready  (slv[3].wready),
      .mst3_wlast   (slv[3].wlast),
      .mst3_wdata   (slv[3].wdata),
      .mst3_wstrb   (slv[3].wstrb),
      .mst3_wuser   (slv[3].wuser),
      .mst3_bvalid  (slv[3].bvalid),
      .mst3_bready  (slv[3].bready),
      .mst3_bid     (slv[3].bid),
      .mst3_bresp   (slv[3].bresp),
      .mst3_buser   (slv[3].buser),
      .mst3_arvalid (slv[3].arvalid),
      .mst3_arready (slv[3].arready),
      .mst3_araddr  (slv[3].araddr),
      .mst3_arlen   (slv[3].arlen),
      .mst3_arsize  (slv[3].arsize),
      .mst3_arburst (slv[3].arburst),
      .mst3_arlock  (slv[3].arlock),
      .mst3_arcache (slv[3].arcache),
      .mst3_arprot  (slv[3].arprot),
      .mst3_arqos   (slv[3].arqos),
      .mst3_arregion(slv[3].arregion),
      .mst3_arid    (slv[3].arid),
      .mst3_aruser  (slv[3].aruser),
      .mst3_rvalid  (slv[3].rvalid),
      .mst3_rready  (slv[3].rready),
      .mst3_rid     (slv[3].rid),
      .mst3_rresp   (slv[3].rresp),
      .mst3_rdata   (slv[3].rdata),
      .mst3_rlast   (slv[3].rlast),
      .mst3_ruser   (slv[3].ruser)
  );

  always #5 aclk = ~aclk;

  initial begin
    aclk = 1'b0;
    aresetn = 1'b1;  // deasserted
    srst = 1'b0;  // deasserted

    // ---For Code Coverage---
    repeat (2) @(posedge aclk);
    srst <= 1'b1;  // asserted
    repeat (10) @(posedge aclk);
    srst <= 1'b0;  // deasserted
    // ---For Code Coverage---

    // Active low reset
    repeat (2) @(posedge aclk);
    aresetn <= 1'b0;  // asserted
    repeat (10) @(posedge aclk);
    aresetn <= 1'b1;  // deasserted
  end

  generate
    for (genvar i = 0; i < 4; i++) begin : gen_config_vif
      initial begin
        uvm_config_db#(virtual axi_if #(AXI_DATA_W, AXI_ADDR_W, AXI_ID_W, AXI_USER_W))::set(
            null, $sformatf("*.master_agent[%0d]", i), "vif", mst[i]);
        uvm_config_db#(virtual axi_if #(AXI_DATA_W, AXI_ADDR_W, AXI_ID_W, AXI_USER_W))::set(
            null, $sformatf("*.slave_agent[%0d]", i), "vif", slv[i]);
      end
    end
  endgenerate

  initial begin
    run_test();
  end


  initial begin
    $fsdbDumpfile("sim.fsdb");
    $fsdbDumpvars();
    $fsdbDumpSVA();
  end

endmodule
