`define DRIVER

class axi_m_driver #(
    int WIDTH = 32,
    SIZE = 3
) extends uvm_driver#(axi_transaction#(WIDTH, SIZE));

  `uvm_component_utils_begin(axi_m_driver#(WIDTH, SIZE))
  `uvm_component_utils_end
  
   axi_subscriber#(WIDTH, SIZE) sub;

  virtual interface axi_intf #(WIDTH, SIZE) intf;

  uvm_analysis_port #(axi_transaction #(WIDTH, SIZE)) drv2sb_port1;
  uvm_analysis_port #(axi_transaction #(WIDTH, SIZE)) drv2sb_port2;


  // new
  int RW;

  axi_transaction #(WIDTH, SIZE) tx;

  function new(string name = "axi_m_driver", uvm_component parent);
    super.new(name, parent);
  endfunction : new

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    drv2sb_port1 = new("drv2sb_port1", this);
    drv2sb_port2 = new("drv2sb_port2", this);
	sub = axi_subscriber#(WIDTH, SIZE)::type_id::create("sub", this);
  endfunction : build_phase


  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    if (!uvm_config_db#(virtual interface axi_intf #(WIDTH, SIZE))::get(this, "", "intf", intf))
      `uvm_error("NOVIF", {"virtual interface must be set for: ", get_full_name(), ".intf"})
	sub.write(intf);
	
  endfunction : connect_phase

  task run_phase(uvm_phase phase);
	super.run_phase(phase);
	// fork
		// reset_intf();
	// join_none
	fork
		sub.do_sample();
		my_send_drv_msg();
	join
  endtask : run_phase
  
  task reset_intf();
	  forever begin
		@(negedge intf.reset) 
  for (int i = 0; i < 3; i++) begin
		intf.M_AWVALID[i] <= 1'b0;
		intf.M_WVALID[i] <= 1'bz;
		intf.M_BREADY[i] = 1'b0;
		intf.M_ARVALID[i] <= 1'b0;
	end
  	end

  endtask

  
  task my_send_drv_msg();
  forever begin
    seq_item_port.get_next_item(req);

/*
    @(posedge intf.clk) 
	  req.RDATA = req.WDATA;
    req.ARADDR = req.AWADDR;
    req.ARLEN = req.AWLEN;
    req.ARSIZE = req.AWSIZE;
    req.ARBURST = req.AWBURST;
*/
    $display("drv seq print:");
    req.print();

	begin 

      sent_addr_write_trx();
      sent_addr_read_trx();
      clr_addr_trx();
      send_data();
     // clr_data();
      send_bresp();
    // clr_bresp();
    //  drv2sb_port1.write(req);
  end

	seq_item_port.item_done();
   	seq_item_port.put(req);
  end
  endtask

  task sent_trx_to_seq();
    begin
      case (RW)
        0: drv2sb_port1.write(req); //RW=0,写操作
        1: drv2sb_port2.write(req); //RW=1,读操作
      endcase
    end
  endtask

//发送写地址
task sent_addr_write_trx();

if(req.M_AWVALID[0])begin  //发送M0写地址到DUT
  		@(posedge intf.clk) begin

			intf.M_AWVALID[0] <= req.M_AWVALID[0];
			intf.M_AWADDR[0] <= req.M_AWADDR[0];
			intf.M_AWBURST[0] <= req.M_AWBURST[0];
			intf.M_AWSIZE[0] <= req.M_AWSIZE[0];                                                             
			intf.M_AWLEN[0] <= req.M_AWLEN[0];
			intf.M_AWID[0] <= req.M_AWID[0];
	end
end

if(req.M_AWVALID[1])begin  //发送M1写地址到DUT
  		@(posedge intf.clk) begin

			intf.M_AWVALID[1] <= req.M_AWVALID[1];
			intf.M_AWADDR[1] <= req.M_AWADDR[1];
			intf.M_AWBURST[1] <= req.M_AWBURST[1];
			intf.M_AWSIZE[1] <= req.M_AWSIZE[1];                                                             
			intf.M_AWLEN[1] <= req.M_AWLEN[1];
			intf.M_AWID[1] <= req.M_AWID[1];
	end
end

if(req.M_AWVALID[2])begin  //发送M2写地址到DUT
  		@(posedge intf.clk) begin

			intf.M_AWVALID[2] <= req.M_AWVALID[2];
			intf.M_AWADDR[2] <= req.M_AWADDR[2];
			intf.M_AWBURST[2] <= req.M_AWBURST[2];
			intf.M_AWSIZE[2] <= req.M_AWSIZE[2];                                                             
			intf.M_AWLEN[2] <= req.M_AWLEN[2];
			intf.M_AWID[2] <= req.M_AWID[2];
	end
end  

  endtask


//发送读地址
  task sent_addr_read_trx();  //发送读地址到DUT

  if(req.M_ARVALID[0])begin  //发送M0读地址到DUT
    @(posedge intf.clk) begin

	    intf.M_ARVALID[0] <= req.M_ARVALID[0];
      intf.M_ARADDR[0] <= req.M_ARADDR[0];
      intf.M_ARLEN[0] <= req.M_ARLEN[0];
	    intf.M_ARBURST[0] <= req.M_ARBURST[0];
      intf.M_ARSIZE[0] <= req.M_ARSIZE[0];
      intf.M_ARID[0] <= req.M_ARID[0];
  end   
    end

  if(req.M_ARVALID[1])begin  //发送M1读地址到DUT
    @(posedge intf.clk) begin

	    intf.M_ARVALID[1] <= req.M_ARVALID[1];
      intf.M_ARADDR[1] <= req.M_ARADDR[1];
      intf.M_ARLEN[1] <= req.M_ARLEN[1];
	    intf.M_ARBURST[1] <= req.M_ARBURST[1];
      intf.M_ARSIZE[1] <= req.M_ARSIZE[1];
      intf.M_ARID[1] <= req.M_ARID[1];
  end   
    end

  if(req.M_ARVALID[2])begin  //发送M2读地址到DUT
    @(posedge intf.clk) begin

	    intf.M_ARVALID[2] <= req.M_ARVALID[2];
      intf.M_ARADDR[2] <= req.M_ARADDR[2];
      intf.M_ARLEN[2] <= req.M_ARLEN[2];
	    intf.M_ARBURST[2] <= req.M_ARBURST[2];
      intf.M_ARSIZE[2] <= req.M_ARSIZE[2];
      intf.M_ARID[2] <= req.M_ARID[2];
  end   
    end

  endtask
  
//清除地址
task clr_addr_trx();

//清除写地址
 
			 @(posedge intf.clk ) 
      if(intf.M_AWREADY[0]) begin 
  
			intf.M_AWVALID[0] <= 'd0;
			intf.M_AWBURST[0] <= 'd0;
			intf.M_AWSIZE[0] <= 'd0;
			intf.M_AWLEN[0] <= 'd0;
			intf.M_AWID[0] <= 'd0;
			intf.M_AWADDR[0] <= 'd0;
			$display("sent addr m0 done");
	end

       if (intf.M_AWREADY[1]) begin
			intf.M_AWVALID[1] <= 'd0;
			intf.M_AWBURST[1] <= 'd0;
			intf.M_AWSIZE[1] <= 'd0;
			intf.M_AWLEN[1] <= 'd0;
			intf.M_AWID[1] <= 'd0;
			intf.M_AWADDR[1] <= 'd0;
			$display("sent addr m1 done");
	end

 
     if (intf.M_AWREADY[2]) begin
			intf.M_AWVALID[2] <= 'd0;
			intf.M_AWBURST[2] <= 'd0;
			intf.M_AWSIZE[2] <= 'd0;
			intf.M_AWLEN[2] <= 'd0;
			intf.M_AWID[2] <= 'd0;
			intf.M_AWADDR[2] <= 'd0;
			$display("sent addr m2 done");
	end

//清除读地址

    if (intf.M_ARREADY[0]) begin
	    intf.M_ARVALID[0] <= 'd0;
      intf.M_ARADDR[0] <= 'd0;
      intf.M_ARLEN[0] <= 'd0;
      intf.M_ARBURST[0] <= 'd0;
      intf.M_ARSIZE[0] <= 'd0;
      intf.M_ARID[0] <= 'd0;
      $display("sent addr m0 read done");
  end   

    if (intf.M_ARREADY[1]) begin
	    intf.M_ARVALID[1] <= 'd0;
      intf.M_ARADDR[1] <= 'd0;
      intf.M_ARLEN[1] <= 'd0;
      intf.M_ARBURST[1] <= 'd0;
      intf.M_ARSIZE[1] <= 'd0;
      intf.M_ARID[1] <= 'd0;
      $display("sent addr m1 read done");
  end   
  
 
     if (intf.M_ARREADY[2])  begin
	    intf.M_ARVALID[2] <= 'd0;
      intf.M_ARADDR[2] <= 'd0;
      intf.M_ARLEN[2] <= 'd0;
      intf.M_ARBURST[2] <= 'd0;
      intf.M_ARSIZE[2] <= 'd0;
      intf.M_ARID[2] <= 'd0;
      $display("sent addr m2 read done");
  end   
endtask


task send_data();

	  if(req.M_WVALID[0] == 1)begin//驱动m0写数据
	    $display("write data m0 start");
      @(posedge intf.clk) 
      begin
        intf.M_WVALID[0] <= req.M_WVALID[0];
        intf.M_WSTRB[0] <= req.M_WSTRB[0];//选中哪几个字写入
        intf.M_WID[0] <= req.M_WID[0];
        intf.M_WDATA[0] <= req.M_WDATA[0];
        intf.M_WLAST[0] <= req.M_WLAST[0];
    end
     end

	  if(req.M_WVALID[1] == 1)begin//驱动m1写数据
	    $display("write data m1 start");
      @(posedge intf.clk)
      begin
        intf.M_WVALID[1] <= req.M_WVALID[1];
        intf.M_WSTRB[1] <= req.M_WSTRB[1];//选中哪几个字写入
        intf.M_WID[1] <= req.M_WID[1];
        intf.M_WDATA[1] <= req.M_WDATA[1];
        intf.M_WLAST[1] <= req.M_WLAST[1];
      end
       end

	  if(req.M_WVALID[2] == 1)begin//驱动m2写数据
	    $display("write data m1 start");
      @(posedge intf.clk) 
      begin
        intf.M_WVALID[2] <= req.M_WVALID[2];
        intf.M_WSTRB[2] <= req.M_WSTRB[2];//选中哪几个字写入
        intf.M_WID[2] <= req.M_WID[2];
        intf.M_WDATA[2] <= req.M_WDATA[2];
        intf.M_WLAST[2] <= req.M_WLAST[2];
      end
         end

//发送读数据
    if(req.S_RVALID[0] == 1 )begin //驱动s0读数据
    $display("read s0 data start");
    @(posedge intf.clk) 
    begin
      intf.S_RVALID[0] <= req.S_RVALID[0];
      intf.S_RID[0]    <= req.S_RID[0];
      intf.S_RDATA[0]  <= req.S_RDATA[0];
      intf.S_RRESP[0]  <= req.S_RRESP[0];
      intf.S_RLAST[0]  <= req.S_RLAST[0];
	  end    
     end

    if(req.S_RVALID[2] == 1 )begin //驱动s2读数据
    $display("read s2 data start");
    @(posedge intf.clk) 
    begin
      intf.S_RVALID[2] <= req.S_RVALID[2];
      intf.S_RID[2]    <= req.S_RID[2];
      intf.S_RDATA[2]  <= req.S_RDATA[2];
      intf.S_RRESP[2]  <= req.S_RRESP[2];
      intf.S_RLAST[2]  <= req.S_RLAST[2];
    end
     end
endtask

//清除数据
task clr_data();

//清除写数据
    begin
        @(posedge intf.clk iff (intf.M_WREADY[0]))
   
        intf.M_WVALID[0] <= 'b0;
        intf.M_WSTRB[0] <= 'b0;
        intf.M_WID[0] <= 'b0;
        intf.M_WDATA[0] <= 'b0;
        intf.M_WLAST[0] <= 'b0;
        $display("write data m0 done");
    end
    begin
        @(posedge intf.clk iff (intf.M_WREADY[1]))
    
        intf.M_WVALID[1] <= 'b0;
        intf.M_WSTRB[1] <= 'b0;
        intf.M_WID[1] <= 'b0;
        intf.M_WDATA[1] <= 'b0;
        intf.M_WLAST[1] <= 'b0;
        $display("write data m1 done");
    end    
    begin
        @(posedge intf.clk iff (intf.M_WREADY[2]))
    
        intf.M_WVALID[2] <= 'b0;
        intf.M_WSTRB[2] <= 'b0;
        intf.M_WID[2] <= 'b0;
        intf.M_WDATA[2] <= 'b0;
        intf.M_WLAST[2] <= 'b0;
        $display("write data m2 done");
    end    

//清除读数据
    begin  
	   @(posedge intf.clk iff (intf.S_RREADY[0]) )
    
      intf.S_RVALID[0] <= 'b0;
      intf.S_RID[0] <= 'b0;
      intf.S_RDATA[0] <= 'b0;
      intf.S_RRESP[0] <= 'b0;
      intf.S_RLAST[0] <= 'b0;
	  $display("read s0 data done");
	  end    

	   @(posedge intf.clk iff (intf.S_RREADY[1]) )
    begin
      intf.S_RVALID[1] <= 'b0;
      intf.S_RID[1] <= 'b0;
      intf.S_RDATA[1] <= 'b0;
      intf.S_RRESP[1] <= 'b0;
      intf.S_RLAST[1] <= 'b0;
    end 

	   @(posedge intf.clk iff (intf.S_RREADY[2]) )
    begin
      intf.S_RVALID[2] <= 'b0;
      intf.S_RID[2] <= 'b0;
      intf.S_RDATA[2] <= 'b0;
      intf.S_RRESP[2] <= 'b0;
      intf.S_RLAST[2] <= 'b0;
	  end    

endtask


task send_bresp();  //发送写响应

		  if(req.S_BVALID[0] == 1'b1) begin
        $display("received write m0 resp start");
        while (!(intf.S_WLAST[0] & intf.S_WREADY[0] & intf.S_WVALID[0])) @(posedge intf.clk);
        intf.S_BID[0] <= req.S_BID[0];
        intf.S_BVALID[0] <= req.S_BVALID[0];
        intf.S_BRESP[0] <= req.S_BRESP[0];
        drv2sb_port1.write(req);//传递m0写响应
        $display("received write m0 resp done");
      end

		  if(req.S_BVALID[1] == 1'b1) begin
        $display("received write m1 resp start");
        while (!(intf.S_WLAST[1] & intf.S_WREADY[1] & intf.S_WVALID[1])) @(posedge intf.clk);
        intf.S_BID[1] <= req.S_BID[1];
        intf.S_BVALID[1] <= req.S_BVALID[1];
        intf.S_BRESP[1] <= req.S_BRESP[1];
        drv2sb_port1.write(req);//传递m1写响应
        $display("received write m1 resp done");
      end

		  if(req.S_BVALID[2] == 1'b1) begin
        $display("received write m2 resp start");
        while (!(intf.S_WLAST[2] & intf.S_WREADY[2] & intf.S_WVALID[2])) @(posedge intf.clk);
        intf.S_BID[2] <= req.S_BID[2];
        intf.S_BVALID[2] <= req.S_BVALID[2];
        intf.S_BRESP[2] <= req.S_BRESP[2];
        drv2sb_port1.write(req);//传递m2写响应
        $display("received write m2 resp done");
      end

endtask

//清除响应
task clr_bresp();

       @(posedge intf.clk iff (intf.S_BVALID[0]))
      begin
        intf.S_BID[0] <= 0;
        intf.S_BVALID[0] <= 0;
        intf.S_BRESP[0] <= 0;	
        $display("received m0 write resp done");
      end
  
       @(posedge intf.clk iff (intf.S_BVALID[1])) 
      begin
        intf.S_BID[1] <= 0;
        intf.S_BVALID[1] <= 0;
        intf.S_BRESP[1] <= 0;	
        $display("received m1 write resp done");
      end

       @(posedge intf.clk iff (intf.S_BVALID[2])) 
      begin
        intf.S_BID[2] <= 0;
        intf.S_BVALID[2] <= 0;
        intf.S_BRESP[2] <= 0;	
       $display("received m2 write resp done");
      end

endtask


endclass

