
`define WIDTH 32 
`define SIZE 3






